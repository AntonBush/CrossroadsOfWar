DADCABABACCBADAAADAAADADRRACBAACABDCACDAACDBADBDBAACACDBADBDBAACADDBADADADCBADBCBAACADBDACBBADCCACCBBAACACCDACBBADABACCBBAAABAACABCBADAAACCBACBBADBDACCBBAACACCAADADADACADCABAACADABADADADCCACCBBAACADBDADADADABACCBADCAACDAACDBADACACCDBAACACBDDADBADDD
ABABADADADCBADBCADBDDADBBAACAABA
ABBCACDBADACADCBADCAACCBADBDDADBBAACAAADAAAC
AADCACBBADDBADBDDADBBAACAAAB
DADCABCBADAAACBBADDBACCBADBCADDD
ABCBADAAACBBADDBACCBADBCAACCACDAACCBACBBADAAADCAACDADADBBAACAABCAACB
ABCBADAAACBBADDBACCBADBCAACCADDADADBBAACBAABAAABAAACBAAAAACAAAAAAABCAAACAAAC
ABCBADAAACBBADDBACCBADBCAACCADDBDADBBAACBAABAAAABAAAAACBAABDAACBAACBAACBAACBAABB
ABCBADAAACBBADDBACCBADBCAACCADDCDADBBAACAAAA
ABCBADAAACBBADDBACCBADBCAACCADABACBBADBCACCBDADBBAACAAAA
ABCBADAAACBBADDBACCBADBCAACCACBCACCBACBBADBCACCADADBBAACAAAA
ABCBADAAACBBADDBACCBADBCAACCACDAACBBACDBADBCDADBBAACAAAA
ABCBADAAACBBADDBACCBADBCAACCACDAACBBACDBADBCAADBADADADAAADADADBCAACCADBCACCBACCADADBBAACAAAABAAAAAABAAAAAAAAAABBAABDAAACAABA
ABCBADAAACBBADDBACCBADBCAACCACDAACBBACDBADBCAADBADADADAAADADADBCAACCACCDADBCACCBACCBADACDADBBAACAAAABAAAAABBAAAAAABCAAACAACBAAACAABA
ABCBADAAACBBADDBACCBADBCAACCACDAACBBACDBADBCAADBADADADAAADADADBCAACCACBCADAAADCBACCBDADBBAACAAAABAAAAAABAACBAACBAAABAABAAAAAAACA
ABCBADAAACBBADDBACCBADBCAACCACBCADADACCAADDBAADBADADADAAADADADBCAACCADBCACCBACCADADBBAACAAAABAAAAABBAABCAABCAABBAABAAAACAABD
ABCBADAAACBBADDBACCBADBCAACCACBCADADACCAADDBAADBADADADAAADADADBCAACCACCDADBCACCBACCBADACDADBBAACAAAABAAAAAADAABCAABAAAADAABDAABAAACA
ABCBADAAACBBADDBACCBADBCAACCACBCADADACCAADDBAADBADADADAAADADADBCAACCACBCADAAADCBACCBDADBBAACAAAABAAAAABDAAAAAAAAAABBAAABAACB
ABCBADAAACBBADDBACCBADBCAACCACCCADAAACBBACCDAADBADADADAAADADADBCAACCADBCACCBACCADADBBAACAAAABAAAAABBAACAAAACAAABAAAAAAACAABC
ABCBADAAACBBADDBACCBADBCAACCACCCADAAACBBACCDAADBADADADAAADADADBCAACCACCDADBCACCBACCBADACDADBBAACAAAABAAAAAAAAABBAABAAAACAAADAABAAAABAABB
ABCBADAAACBBADDBACCBADBCAACCACCCADAAACBBACCDAADBADADADAAADADADBCAACCACBCADAAADCBACCBDADBBAACAAAABAAAAABDAABCAACBAAADAABBAACBAABB
ABCBADAAACBBADDBACCBADBCAACCACCBADDBACCBADBDAADBADADADAAADADADBCAACCADBCACCBACCADADBBAACAAAABAAAAABCAAACAAACAACAAABBAABBAABC
ABCBADAAACBBADDBACCBADBCAACCACCBADDBACCBADBDAADBADADADAAADADADBCAACCACCDADBCACCBACCBADACDADBBAACAAAABAAAAACAAABBAACAAABAAAACAABBAABC
ABCBADAAACBBADDBACCBADBCAACCACCBADDBACCBADBDAADBADADADAAADADADBCAACCACBCADAAADCBACCBDADBBAACAAAABAAAAABCAAAAAACBAACBAABDAABBAACB
ABCBADAAACBBADDBACCBADBCAACCACDAACBBADBDAADAADADADCDDADBBAACAAAA
ABCBADADADACACDBACCBADBDAADBADADADCBADACADCADADBBAACAAAA
ABABADCBADACADCAACCBADBCADBDAADBADADADCBADACADCADADBBAACAAAA
DADCABCAADCAACDAACCBADBCAADBADBCACCBACBBADCAADCBADBCACCBADBDADDD
ABDDADACACDBABDBADBAACBBADCDADACAACCACDAACCBACBBADAAADCAACDADADBBAACAACAAAAAAAAA
ABDCACDBADABACBCACCBADBCAAABAACCACDAACCBACBBADAAADCAACDADADBBAACAAABAABCAAAA
ABDCACDBADABACBCACCBADBCAAACAACCACDAACCBACBBADAAADCAACDADADBBAACAAABAABCAAAA
ABDDADBCADBDACBBAACCACDAACCBACBBADAAADCAACDADADBBAACAAACAAAAAAAAAAAA
DADCABDAACCBADBDADADADCBADBCADBDACCBADBDADDD
ACABADADADADACCADADBBAACAAAA
DDAAADADADADACCADADBBAACAAAA
DADCABACADCAACCBADABADBDADDD
ABACADCAACCBADABADBDAADBADADADCBADACADCADADBBAACAAAA
DADCAADAADCBACDBADAAACCAACDBADACACCDADBDADDD
DDAAACDBADBCACCBABBBACCBADCCACCBADAADADBBAACAAAB
ACABACBBADBCACCBACDAADADADCBADBDACCBDADBBAACAAAA
ACABACCBACBBADBAADADADACDADBBAACAAAA
DDAAACBBADBCADABDADBBAACAAAA
ABABADADADCBADBDACCBADBDDADBBAACAAAA
ABBBACCBACCCADCAABDCADADADCDACCBADBCDADBBAACAAAA
ABDAACDBACCDACDAADCAABDCADADADCDACCBADBCDADBBAACAAAA
ABBBACCBACCCADCAACABACBBADAAADAADADBBAACAAAA
ABBBACCBACCCADCAACABACBBADAAADAAAACCACDAACCBACBBADAAADCAACDADADBBAACAAAA
ABDAACDBACCDACDAADCAACABACBBADAAADAADADBBAACAAAA
ABDAACDBACCDACDAADCAACABACBBADAAADAAAACCACDAACCBACBBADAAADCAACDADADBBAACAAAA
ABDCADBCACCBACCBAACCAAAADADBBAACAAAB
ABDCADBCACCBACCBAACCAAABDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACDADBBAACAAAB
ABDCADBCACCBACCBAACCAAADDADBBAACAAAB
ABDCADBCACCBACCBAACCAABADADBBAACAAAB
ABDCADBCACCBACCBAACCAABBDADBBAACAAAB
ABDCADBCACCBACCBAACCAABCDADBBAACAAAB
ABDCADBCACCBACCBAACCAABDDADBBAACAAAB
ABDCADBCACCBACCBAACCAACADADBBAACAAAB
ABDCADBCACCBACCBAACCAACBDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAAAADADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAAABDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAAACDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAAADDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAABADADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAABBDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAABCDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAABDDADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAACADADBBAACAAAB
ABDCADBCACCBACCBAACCAAABAACBDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAAAADADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAAABDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAAACDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAAADDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAABADADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAABBDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAABCDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAABDDADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAACADADBBAACAAAB
ABDCADBCACCBACCBAACCAAACAACBDADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAAAADADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAAABDADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAAACDADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAAADDADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAABADADBBAACAAAB
ABDCADBCACCBACCBAACCAAADAABBDADBBAACAAAB
ADCDACCBACBBADCAACDAACCBADBCDADBBAACAAAA
ABDBADCBADACAACCADDADADBBAACBAABAAACAABCBAAAAAABAABAAABAAACAAABC
ABDBADCBADACAACCADDBDADBBAACAAACBAAAAAABAABAAABDAABDAABDAAAD
DADCABBCADCBADBDACDBACBDADDD
ABBCADCBADBDACDBACBDAACCABBBADCCADADDADBBAACAAAA
ABBCADCBADBDACDBACBDAACCABBBADCCAAACDADBBAACAAAA
ABBCADCBADBDACDBACBDAACCABBBADCCAAADDADBBAACAAAA
ABBCADCBADBDACDBACBDAACCDDAAACDBACCDACDAADCADADBBAACAAAA
ABBCADCBADBDACDBACBDAACCABDBACBBACCADADBBAACAAAA
